`include "define.v"

module ID(
	
);