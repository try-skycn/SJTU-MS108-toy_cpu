module MIPS(
	input	wire	clk,
	input	wire	rst
);

/*
	compile module CPU
	compile module InstRom
	compile module DataRam
*/

endmodule
